module FullAdder(a,b,cin,cout,sum);
endmodule